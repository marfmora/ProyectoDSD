-- Sistema_Epy.vhd

-- Generated using ACDS version 16.1 196

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Sistema_Epy is
	port (
		clk_clk                      : in    std_logic                     := '0';             --                    clk.clk
		clk_sdram_clk                : out   std_logic;                                        --              clk_sdram.clk
		reset_reset_n                : in    std_logic                     := '0';             --                  reset.reset_n
		sdram_wire_addr              : out   std_logic_vector(12 downto 0);                    --             sdram_wire.addr
		sdram_wire_ba                : out   std_logic_vector(1 downto 0);                     --                       .ba
		sdram_wire_cas_n             : out   std_logic;                                        --                       .cas_n
		sdram_wire_cke               : out   std_logic;                                        --                       .cke
		sdram_wire_cs_n              : out   std_logic;                                        --                       .cs_n
		sdram_wire_dq                : inout std_logic_vector(15 downto 0) := (others => '0'); --                       .dq
		sdram_wire_dqm               : out   std_logic_vector(1 downto 0);                     --                       .dqm
		sdram_wire_ras_n             : out   std_logic;                                        --                       .ras_n
		sdram_wire_we_n              : out   std_logic;                                        --                       .we_n
		uart_rxd                     : in    std_logic                     := '0';             --                   uart.rxd
		uart_txd                     : out   std_logic;                                        --                       .txd
		vga_external_interface_CLK   : out   std_logic;                                        -- vga_external_interface.CLK
		vga_external_interface_HS    : out   std_logic;                                        --                       .HS
		vga_external_interface_VS    : out   std_logic;                                        --                       .VS
		vga_external_interface_BLANK : out   std_logic;                                        --                       .BLANK
		vga_external_interface_SYNC  : out   std_logic;                                        --                       .SYNC
		vga_external_interface_R     : out   std_logic_vector(7 downto 0);                     --                       .R
		vga_external_interface_G     : out   std_logic_vector(7 downto 0);                     --                       .G
		vga_external_interface_B     : out   std_logic_vector(7 downto 0)                      --                       .B
	);
end entity Sistema_Epy;

architecture rtl of Sistema_Epy is
	component Sistema_Epy_DUAL_CLOCK_FIFO is
		port (
			clk_stream_in            : in  std_logic                     := 'X';             -- clk
			reset_stream_in          : in  std_logic                     := 'X';             -- reset
			clk_stream_out           : in  std_logic                     := 'X';             -- clk
			reset_stream_out         : in  std_logic                     := 'X';             -- reset
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_data           : in  std_logic_vector(29 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(29 downto 0)                     -- data
		);
	end component Sistema_Epy_DUAL_CLOCK_FIFO;

	component Sistema_Epy_JTAG_UART is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component Sistema_Epy_JTAG_UART;

	component Sistema_Epy_NIOS2_NN is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(19 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(19 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component Sistema_Epy_NIOS2_NN;

	component Sistema_Epy_NIOS2_VGA is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(26 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(19 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component Sistema_Epy_NIOS2_VGA;

	component Sistema_Epy_PIXEL_BUFFER_DMA is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_arbiterlock   : out std_logic;                                        -- lock
			master_read          : out std_logic;                                        -- read
			master_readdata      : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			slave_address        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			slave_byteenable     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			slave_read           : in  std_logic                     := 'X';             -- read
			slave_write          : in  std_logic                     := 'X';             -- write
			slave_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			slave_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			stream_ready         : in  std_logic                     := 'X';             -- ready
			stream_startofpacket : out std_logic;                                        -- startofpacket
			stream_endofpacket   : out std_logic;                                        -- endofpacket
			stream_valid         : out std_logic;                                        -- valid
			stream_data          : out std_logic_vector(15 downto 0)                     -- data
		);
	end component Sistema_Epy_PIXEL_BUFFER_DMA;

	component Sistema_Epy_PLL is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			outclk_1 : out std_logic;        -- clk
			outclk_2 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component Sistema_Epy_PLL;

	component Sistema_Epy_RGB_RESAMPLER is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_data           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(29 downto 0)                     -- data
		);
	end component Sistema_Epy_RGB_RESAMPLER;

	component Sistema_Epy_SCALER is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_data           : in  std_logic_vector(29 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(29 downto 0);                    -- data
			stream_out_channel       : out std_logic_vector(1 downto 0)                      -- channel
		);
	end component Sistema_Epy_SCALER;

	component Sistema_Epy_SDRAM_VGA is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component Sistema_Epy_SDRAM_VGA;

	component Sistema_Epy_SYSTEM_ID_1 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component Sistema_Epy_SYSTEM_ID_1;

	component Sistema_Epy_TIMER is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component Sistema_Epy_TIMER;

	component Sistema_Epy_VGA is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset         : in  std_logic                     := 'X';             -- reset
			data          : in  std_logic_vector(29 downto 0) := (others => 'X'); -- data
			startofpacket : in  std_logic                     := 'X';             -- startofpacket
			endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			valid         : in  std_logic                     := 'X';             -- valid
			ready         : out std_logic;                                        -- ready
			VGA_CLK       : out std_logic;                                        -- export
			VGA_HS        : out std_logic;                                        -- export
			VGA_VS        : out std_logic;                                        -- export
			VGA_BLANK     : out std_logic;                                        -- export
			VGA_SYNC      : out std_logic;                                        -- export
			VGA_R         : out std_logic_vector(7 downto 0);                     -- export
			VGA_G         : out std_logic_vector(7 downto 0);                     -- export
			VGA_B         : out std_logic_vector(7 downto 0)                      -- export
		);
	end component Sistema_Epy_VGA;

	component Sistema_Epy_onchip_mem2 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component Sistema_Epy_onchip_mem2;

	component Sistema_Epy_onchip_mem3 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component Sistema_Epy_onchip_mem3;

	component Sistema_Epy_uart_0 is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			read_n        : in  std_logic                     := 'X';             -- read_n
			write_n       : in  std_logic                     := 'X';             -- write_n
			writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			rxd           : in  std_logic                     := 'X';             -- export
			txd           : out std_logic;                                        -- export
			irq           : out std_logic                                         -- irq
		);
	end component Sistema_Epy_uart_0;

	component Sistema_Epy_mm_interconnect_0 is
		port (
			PLL_outclk0_clk                                        : in  std_logic                     := 'X';             -- clk
			PIXEL_BUFFER_DMA_reset_reset_bridge_in_reset_reset     : in  std_logic                     := 'X';             -- reset
			NIOS2_NN_data_master_address                           : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			NIOS2_NN_data_master_waitrequest                       : out std_logic;                                        -- waitrequest
			NIOS2_NN_data_master_byteenable                        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			NIOS2_NN_data_master_read                              : in  std_logic                     := 'X';             -- read
			NIOS2_NN_data_master_readdata                          : out std_logic_vector(31 downto 0);                    -- readdata
			NIOS2_NN_data_master_write                             : in  std_logic                     := 'X';             -- write
			NIOS2_NN_data_master_writedata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			NIOS2_NN_data_master_debugaccess                       : in  std_logic                     := 'X';             -- debugaccess
			NIOS2_NN_instruction_master_address                    : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			NIOS2_NN_instruction_master_waitrequest                : out std_logic;                                        -- waitrequest
			NIOS2_NN_instruction_master_read                       : in  std_logic                     := 'X';             -- read
			NIOS2_NN_instruction_master_readdata                   : out std_logic_vector(31 downto 0);                    -- readdata
			NIOS2_VGA_data_master_address                          : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			NIOS2_VGA_data_master_waitrequest                      : out std_logic;                                        -- waitrequest
			NIOS2_VGA_data_master_byteenable                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			NIOS2_VGA_data_master_read                             : in  std_logic                     := 'X';             -- read
			NIOS2_VGA_data_master_readdata                         : out std_logic_vector(31 downto 0);                    -- readdata
			NIOS2_VGA_data_master_readdatavalid                    : out std_logic;                                        -- readdatavalid
			NIOS2_VGA_data_master_write                            : in  std_logic                     := 'X';             -- write
			NIOS2_VGA_data_master_writedata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			NIOS2_VGA_data_master_debugaccess                      : in  std_logic                     := 'X';             -- debugaccess
			NIOS2_VGA_instruction_master_address                   : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			NIOS2_VGA_instruction_master_waitrequest               : out std_logic;                                        -- waitrequest
			NIOS2_VGA_instruction_master_read                      : in  std_logic                     := 'X';             -- read
			NIOS2_VGA_instruction_master_readdata                  : out std_logic_vector(31 downto 0);                    -- readdata
			NIOS2_VGA_instruction_master_readdatavalid             : out std_logic;                                        -- readdatavalid
			PIXEL_BUFFER_DMA_avalon_pixel_dma_master_address       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			PIXEL_BUFFER_DMA_avalon_pixel_dma_master_waitrequest   : out std_logic;                                        -- waitrequest
			PIXEL_BUFFER_DMA_avalon_pixel_dma_master_read          : in  std_logic                     := 'X';             -- read
			PIXEL_BUFFER_DMA_avalon_pixel_dma_master_readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			PIXEL_BUFFER_DMA_avalon_pixel_dma_master_readdatavalid : out std_logic;                                        -- readdatavalid
			PIXEL_BUFFER_DMA_avalon_pixel_dma_master_lock          : in  std_logic                     := 'X';             -- lock
			JTAG_UART_avalon_jtag_slave_address                    : out std_logic_vector(0 downto 0);                     -- address
			JTAG_UART_avalon_jtag_slave_write                      : out std_logic;                                        -- write
			JTAG_UART_avalon_jtag_slave_read                       : out std_logic;                                        -- read
			JTAG_UART_avalon_jtag_slave_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			JTAG_UART_avalon_jtag_slave_writedata                  : out std_logic_vector(31 downto 0);                    -- writedata
			JTAG_UART_avalon_jtag_slave_waitrequest                : in  std_logic                     := 'X';             -- waitrequest
			JTAG_UART_avalon_jtag_slave_chipselect                 : out std_logic;                                        -- chipselect
			NIOS2_NN_debug_mem_slave_address                       : out std_logic_vector(8 downto 0);                     -- address
			NIOS2_NN_debug_mem_slave_write                         : out std_logic;                                        -- write
			NIOS2_NN_debug_mem_slave_read                          : out std_logic;                                        -- read
			NIOS2_NN_debug_mem_slave_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			NIOS2_NN_debug_mem_slave_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			NIOS2_NN_debug_mem_slave_byteenable                    : out std_logic_vector(3 downto 0);                     -- byteenable
			NIOS2_NN_debug_mem_slave_waitrequest                   : in  std_logic                     := 'X';             -- waitrequest
			NIOS2_NN_debug_mem_slave_debugaccess                   : out std_logic;                                        -- debugaccess
			NIOS2_VGA_debug_mem_slave_address                      : out std_logic_vector(8 downto 0);                     -- address
			NIOS2_VGA_debug_mem_slave_write                        : out std_logic;                                        -- write
			NIOS2_VGA_debug_mem_slave_read                         : out std_logic;                                        -- read
			NIOS2_VGA_debug_mem_slave_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			NIOS2_VGA_debug_mem_slave_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			NIOS2_VGA_debug_mem_slave_byteenable                   : out std_logic_vector(3 downto 0);                     -- byteenable
			NIOS2_VGA_debug_mem_slave_waitrequest                  : in  std_logic                     := 'X';             -- waitrequest
			NIOS2_VGA_debug_mem_slave_debugaccess                  : out std_logic;                                        -- debugaccess
			onchip_mem2_s1_address                                 : out std_logic_vector(15 downto 0);                    -- address
			onchip_mem2_s1_write                                   : out std_logic;                                        -- write
			onchip_mem2_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_mem2_s1_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_mem2_s1_byteenable                              : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_mem2_s1_chipselect                              : out std_logic;                                        -- chipselect
			onchip_mem2_s1_clken                                   : out std_logic;                                        -- clken
			onchip_mem3_s1_address                                 : out std_logic_vector(15 downto 0);                    -- address
			onchip_mem3_s1_write                                   : out std_logic;                                        -- write
			onchip_mem3_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_mem3_s1_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_mem3_s1_byteenable                              : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_mem3_s1_chipselect                              : out std_logic;                                        -- chipselect
			onchip_mem3_s1_clken                                   : out std_logic;                                        -- clken
			PIXEL_BUFFER_DMA_avalon_control_slave_address          : out std_logic_vector(1 downto 0);                     -- address
			PIXEL_BUFFER_DMA_avalon_control_slave_write            : out std_logic;                                        -- write
			PIXEL_BUFFER_DMA_avalon_control_slave_read             : out std_logic;                                        -- read
			PIXEL_BUFFER_DMA_avalon_control_slave_readdata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			PIXEL_BUFFER_DMA_avalon_control_slave_writedata        : out std_logic_vector(31 downto 0);                    -- writedata
			PIXEL_BUFFER_DMA_avalon_control_slave_byteenable       : out std_logic_vector(3 downto 0);                     -- byteenable
			SDRAM_VGA_s1_address                                   : out std_logic_vector(24 downto 0);                    -- address
			SDRAM_VGA_s1_write                                     : out std_logic;                                        -- write
			SDRAM_VGA_s1_read                                      : out std_logic;                                        -- read
			SDRAM_VGA_s1_readdata                                  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			SDRAM_VGA_s1_writedata                                 : out std_logic_vector(15 downto 0);                    -- writedata
			SDRAM_VGA_s1_byteenable                                : out std_logic_vector(1 downto 0);                     -- byteenable
			SDRAM_VGA_s1_readdatavalid                             : in  std_logic                     := 'X';             -- readdatavalid
			SDRAM_VGA_s1_waitrequest                               : in  std_logic                     := 'X';             -- waitrequest
			SDRAM_VGA_s1_chipselect                                : out std_logic;                                        -- chipselect
			SYSTEM_ID_1_control_slave_address                      : out std_logic_vector(0 downto 0);                     -- address
			SYSTEM_ID_1_control_slave_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			TIMER_s1_address                                       : out std_logic_vector(2 downto 0);                     -- address
			TIMER_s1_write                                         : out std_logic;                                        -- write
			TIMER_s1_readdata                                      : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			TIMER_s1_writedata                                     : out std_logic_vector(15 downto 0);                    -- writedata
			TIMER_s1_chipselect                                    : out std_logic                                         -- chipselect
		);
	end component Sistema_Epy_mm_interconnect_0;

	component Sistema_Epy_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component Sistema_Epy_irq_mapper;

	component Sistema_Epy_avalon_st_adapter is
		generic (
			inBitsPerSymbol : integer := 8;
			inUsePackets    : integer := 0;
			inDataWidth     : integer := 8;
			inChannelWidth  : integer := 3;
			inErrorWidth    : integer := 2;
			inUseEmptyPort  : integer := 0;
			inUseValid      : integer := 1;
			inUseReady      : integer := 1;
			inReadyLatency  : integer := 0;
			outDataWidth    : integer := 32;
			outChannelWidth : integer := 3;
			outErrorWidth   : integer := 2;
			outUseEmptyPort : integer := 0;
			outUseValid     : integer := 1;
			outUseReady     : integer := 1;
			outReadyLatency : integer := 0
		);
		port (
			in_clk_0_clk        : in  std_logic                     := 'X';             -- clk
			in_rst_0_reset      : in  std_logic                     := 'X';             -- reset
			in_0_data           : in  std_logic_vector(29 downto 0) := (others => 'X'); -- data
			in_0_valid          : in  std_logic                     := 'X';             -- valid
			in_0_ready          : out std_logic;                                        -- ready
			in_0_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_0_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			in_0_channel        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- channel
			out_0_data          : out std_logic_vector(29 downto 0);                    -- data
			out_0_valid         : out std_logic;                                        -- valid
			out_0_ready         : in  std_logic                     := 'X';             -- ready
			out_0_startofpacket : out std_logic;                                        -- startofpacket
			out_0_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component Sistema_Epy_avalon_st_adapter;

	component sistema_epy_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_in2      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component sistema_epy_rst_controller;

	component sistema_epy_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_in2      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component sistema_epy_rst_controller_001;

	signal dual_clock_fifo_avalon_dc_buffer_source_valid                      : std_logic;                     -- DUAL_CLOCK_FIFO:stream_out_valid -> VGA:valid
	signal dual_clock_fifo_avalon_dc_buffer_source_data                       : std_logic_vector(29 downto 0); -- DUAL_CLOCK_FIFO:stream_out_data -> VGA:data
	signal dual_clock_fifo_avalon_dc_buffer_source_ready                      : std_logic;                     -- VGA:ready -> DUAL_CLOCK_FIFO:stream_out_ready
	signal dual_clock_fifo_avalon_dc_buffer_source_startofpacket              : std_logic;                     -- DUAL_CLOCK_FIFO:stream_out_startofpacket -> VGA:startofpacket
	signal dual_clock_fifo_avalon_dc_buffer_source_endofpacket                : std_logic;                     -- DUAL_CLOCK_FIFO:stream_out_endofpacket -> VGA:endofpacket
	signal pixel_buffer_dma_avalon_pixel_source_valid                         : std_logic;                     -- PIXEL_BUFFER_DMA:stream_valid -> RGB_RESAMPLER:stream_in_valid
	signal pixel_buffer_dma_avalon_pixel_source_data                          : std_logic_vector(15 downto 0); -- PIXEL_BUFFER_DMA:stream_data -> RGB_RESAMPLER:stream_in_data
	signal pixel_buffer_dma_avalon_pixel_source_ready                         : std_logic;                     -- RGB_RESAMPLER:stream_in_ready -> PIXEL_BUFFER_DMA:stream_ready
	signal pixel_buffer_dma_avalon_pixel_source_startofpacket                 : std_logic;                     -- PIXEL_BUFFER_DMA:stream_startofpacket -> RGB_RESAMPLER:stream_in_startofpacket
	signal pixel_buffer_dma_avalon_pixel_source_endofpacket                   : std_logic;                     -- PIXEL_BUFFER_DMA:stream_endofpacket -> RGB_RESAMPLER:stream_in_endofpacket
	signal rgb_resampler_avalon_rgb_source_valid                              : std_logic;                     -- RGB_RESAMPLER:stream_out_valid -> SCALER:stream_in_valid
	signal rgb_resampler_avalon_rgb_source_data                               : std_logic_vector(29 downto 0); -- RGB_RESAMPLER:stream_out_data -> SCALER:stream_in_data
	signal rgb_resampler_avalon_rgb_source_ready                              : std_logic;                     -- SCALER:stream_in_ready -> RGB_RESAMPLER:stream_out_ready
	signal rgb_resampler_avalon_rgb_source_startofpacket                      : std_logic;                     -- RGB_RESAMPLER:stream_out_startofpacket -> SCALER:stream_in_startofpacket
	signal rgb_resampler_avalon_rgb_source_endofpacket                        : std_logic;                     -- RGB_RESAMPLER:stream_out_endofpacket -> SCALER:stream_in_endofpacket
	signal pll_outclk0_clk                                                    : std_logic;                     -- PLL:outclk_0 -> [DUAL_CLOCK_FIFO:clk_stream_in, JTAG_UART:clk, NIOS2_NN:clk, NIOS2_VGA:clk, PIXEL_BUFFER_DMA:clk, RGB_RESAMPLER:clk, SCALER:clk, SDRAM_VGA:clk, SYSTEM_ID_1:clock, TIMER:clk, avalon_st_adapter:in_clk_0_clk, irq_mapper:clk, irq_mapper_001:clk, mm_interconnect_0:PLL_outclk0_clk, onchip_mem2:clk, onchip_mem3:clk, rst_controller:clk, uart_0:clk]
	signal pll_outclk1_clk                                                    : std_logic;                     -- PLL:outclk_1 -> [DUAL_CLOCK_FIFO:clk_stream_out, VGA:clk, rst_controller_001:clk]
	signal pixel_buffer_dma_avalon_pixel_dma_master_waitrequest               : std_logic;                     -- mm_interconnect_0:PIXEL_BUFFER_DMA_avalon_pixel_dma_master_waitrequest -> PIXEL_BUFFER_DMA:master_waitrequest
	signal pixel_buffer_dma_avalon_pixel_dma_master_readdata                  : std_logic_vector(15 downto 0); -- mm_interconnect_0:PIXEL_BUFFER_DMA_avalon_pixel_dma_master_readdata -> PIXEL_BUFFER_DMA:master_readdata
	signal pixel_buffer_dma_avalon_pixel_dma_master_address                   : std_logic_vector(31 downto 0); -- PIXEL_BUFFER_DMA:master_address -> mm_interconnect_0:PIXEL_BUFFER_DMA_avalon_pixel_dma_master_address
	signal pixel_buffer_dma_avalon_pixel_dma_master_read                      : std_logic;                     -- PIXEL_BUFFER_DMA:master_read -> mm_interconnect_0:PIXEL_BUFFER_DMA_avalon_pixel_dma_master_read
	signal pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid             : std_logic;                     -- mm_interconnect_0:PIXEL_BUFFER_DMA_avalon_pixel_dma_master_readdatavalid -> PIXEL_BUFFER_DMA:master_readdatavalid
	signal pixel_buffer_dma_avalon_pixel_dma_master_lock                      : std_logic;                     -- PIXEL_BUFFER_DMA:master_arbiterlock -> mm_interconnect_0:PIXEL_BUFFER_DMA_avalon_pixel_dma_master_lock
	signal nios2_vga_data_master_readdata                                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:NIOS2_VGA_data_master_readdata -> NIOS2_VGA:d_readdata
	signal nios2_vga_data_master_waitrequest                                  : std_logic;                     -- mm_interconnect_0:NIOS2_VGA_data_master_waitrequest -> NIOS2_VGA:d_waitrequest
	signal nios2_vga_data_master_debugaccess                                  : std_logic;                     -- NIOS2_VGA:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NIOS2_VGA_data_master_debugaccess
	signal nios2_vga_data_master_address                                      : std_logic_vector(26 downto 0); -- NIOS2_VGA:d_address -> mm_interconnect_0:NIOS2_VGA_data_master_address
	signal nios2_vga_data_master_byteenable                                   : std_logic_vector(3 downto 0);  -- NIOS2_VGA:d_byteenable -> mm_interconnect_0:NIOS2_VGA_data_master_byteenable
	signal nios2_vga_data_master_read                                         : std_logic;                     -- NIOS2_VGA:d_read -> mm_interconnect_0:NIOS2_VGA_data_master_read
	signal nios2_vga_data_master_readdatavalid                                : std_logic;                     -- mm_interconnect_0:NIOS2_VGA_data_master_readdatavalid -> NIOS2_VGA:d_readdatavalid
	signal nios2_vga_data_master_write                                        : std_logic;                     -- NIOS2_VGA:d_write -> mm_interconnect_0:NIOS2_VGA_data_master_write
	signal nios2_vga_data_master_writedata                                    : std_logic_vector(31 downto 0); -- NIOS2_VGA:d_writedata -> mm_interconnect_0:NIOS2_VGA_data_master_writedata
	signal nios2_nn_data_master_readdata                                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:NIOS2_NN_data_master_readdata -> NIOS2_NN:d_readdata
	signal nios2_nn_data_master_waitrequest                                   : std_logic;                     -- mm_interconnect_0:NIOS2_NN_data_master_waitrequest -> NIOS2_NN:d_waitrequest
	signal nios2_nn_data_master_debugaccess                                   : std_logic;                     -- NIOS2_NN:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NIOS2_NN_data_master_debugaccess
	signal nios2_nn_data_master_address                                       : std_logic_vector(19 downto 0); -- NIOS2_NN:d_address -> mm_interconnect_0:NIOS2_NN_data_master_address
	signal nios2_nn_data_master_byteenable                                    : std_logic_vector(3 downto 0);  -- NIOS2_NN:d_byteenable -> mm_interconnect_0:NIOS2_NN_data_master_byteenable
	signal nios2_nn_data_master_read                                          : std_logic;                     -- NIOS2_NN:d_read -> mm_interconnect_0:NIOS2_NN_data_master_read
	signal nios2_nn_data_master_write                                         : std_logic;                     -- NIOS2_NN:d_write -> mm_interconnect_0:NIOS2_NN_data_master_write
	signal nios2_nn_data_master_writedata                                     : std_logic_vector(31 downto 0); -- NIOS2_NN:d_writedata -> mm_interconnect_0:NIOS2_NN_data_master_writedata
	signal nios2_nn_instruction_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:NIOS2_NN_instruction_master_readdata -> NIOS2_NN:i_readdata
	signal nios2_nn_instruction_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:NIOS2_NN_instruction_master_waitrequest -> NIOS2_NN:i_waitrequest
	signal nios2_nn_instruction_master_address                                : std_logic_vector(19 downto 0); -- NIOS2_NN:i_address -> mm_interconnect_0:NIOS2_NN_instruction_master_address
	signal nios2_nn_instruction_master_read                                   : std_logic;                     -- NIOS2_NN:i_read -> mm_interconnect_0:NIOS2_NN_instruction_master_read
	signal nios2_vga_instruction_master_readdata                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:NIOS2_VGA_instruction_master_readdata -> NIOS2_VGA:i_readdata
	signal nios2_vga_instruction_master_waitrequest                           : std_logic;                     -- mm_interconnect_0:NIOS2_VGA_instruction_master_waitrequest -> NIOS2_VGA:i_waitrequest
	signal nios2_vga_instruction_master_address                               : std_logic_vector(19 downto 0); -- NIOS2_VGA:i_address -> mm_interconnect_0:NIOS2_VGA_instruction_master_address
	signal nios2_vga_instruction_master_read                                  : std_logic;                     -- NIOS2_VGA:i_read -> mm_interconnect_0:NIOS2_VGA_instruction_master_read
	signal nios2_vga_instruction_master_readdatavalid                         : std_logic;                     -- mm_interconnect_0:NIOS2_VGA_instruction_master_readdatavalid -> NIOS2_VGA:i_readdatavalid
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect           : std_logic;                     -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_chipselect -> JTAG_UART:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata             : std_logic_vector(31 downto 0); -- JTAG_UART:av_readdata -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest          : std_logic;                     -- JTAG_UART:av_waitrequest -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address              : std_logic_vector(0 downto 0);  -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_address -> JTAG_UART:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read                 : std_logic;                     -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write                : std_logic;                     -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_writedata -> JTAG_UART:av_writedata
	signal mm_interconnect_0_sdram_vga_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:SDRAM_VGA_s1_chipselect -> SDRAM_VGA:az_cs
	signal mm_interconnect_0_sdram_vga_s1_readdata                            : std_logic_vector(15 downto 0); -- SDRAM_VGA:za_data -> mm_interconnect_0:SDRAM_VGA_s1_readdata
	signal mm_interconnect_0_sdram_vga_s1_waitrequest                         : std_logic;                     -- SDRAM_VGA:za_waitrequest -> mm_interconnect_0:SDRAM_VGA_s1_waitrequest
	signal mm_interconnect_0_sdram_vga_s1_address                             : std_logic_vector(24 downto 0); -- mm_interconnect_0:SDRAM_VGA_s1_address -> SDRAM_VGA:az_addr
	signal mm_interconnect_0_sdram_vga_s1_read                                : std_logic;                     -- mm_interconnect_0:SDRAM_VGA_s1_read -> mm_interconnect_0_sdram_vga_s1_read:in
	signal mm_interconnect_0_sdram_vga_s1_byteenable                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:SDRAM_VGA_s1_byteenable -> mm_interconnect_0_sdram_vga_s1_byteenable:in
	signal mm_interconnect_0_sdram_vga_s1_readdatavalid                       : std_logic;                     -- SDRAM_VGA:za_valid -> mm_interconnect_0:SDRAM_VGA_s1_readdatavalid
	signal mm_interconnect_0_sdram_vga_s1_write                               : std_logic;                     -- mm_interconnect_0:SDRAM_VGA_s1_write -> mm_interconnect_0_sdram_vga_s1_write:in
	signal mm_interconnect_0_sdram_vga_s1_writedata                           : std_logic_vector(15 downto 0); -- mm_interconnect_0:SDRAM_VGA_s1_writedata -> SDRAM_VGA:az_data
	signal mm_interconnect_0_system_id_1_control_slave_readdata               : std_logic_vector(31 downto 0); -- SYSTEM_ID_1:readdata -> mm_interconnect_0:SYSTEM_ID_1_control_slave_readdata
	signal mm_interconnect_0_system_id_1_control_slave_address                : std_logic_vector(0 downto 0);  -- mm_interconnect_0:SYSTEM_ID_1_control_slave_address -> SYSTEM_ID_1:address
	signal mm_interconnect_0_nios2_nn_debug_mem_slave_readdata                : std_logic_vector(31 downto 0); -- NIOS2_NN:debug_mem_slave_readdata -> mm_interconnect_0:NIOS2_NN_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_nn_debug_mem_slave_waitrequest             : std_logic;                     -- NIOS2_NN:debug_mem_slave_waitrequest -> mm_interconnect_0:NIOS2_NN_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_nn_debug_mem_slave_debugaccess             : std_logic;                     -- mm_interconnect_0:NIOS2_NN_debug_mem_slave_debugaccess -> NIOS2_NN:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_nn_debug_mem_slave_address                 : std_logic_vector(8 downto 0);  -- mm_interconnect_0:NIOS2_NN_debug_mem_slave_address -> NIOS2_NN:debug_mem_slave_address
	signal mm_interconnect_0_nios2_nn_debug_mem_slave_read                    : std_logic;                     -- mm_interconnect_0:NIOS2_NN_debug_mem_slave_read -> NIOS2_NN:debug_mem_slave_read
	signal mm_interconnect_0_nios2_nn_debug_mem_slave_byteenable              : std_logic_vector(3 downto 0);  -- mm_interconnect_0:NIOS2_NN_debug_mem_slave_byteenable -> NIOS2_NN:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_nn_debug_mem_slave_write                   : std_logic;                     -- mm_interconnect_0:NIOS2_NN_debug_mem_slave_write -> NIOS2_NN:debug_mem_slave_write
	signal mm_interconnect_0_nios2_nn_debug_mem_slave_writedata               : std_logic_vector(31 downto 0); -- mm_interconnect_0:NIOS2_NN_debug_mem_slave_writedata -> NIOS2_NN:debug_mem_slave_writedata
	signal mm_interconnect_0_timer_s1_chipselect                              : std_logic;                     -- mm_interconnect_0:TIMER_s1_chipselect -> TIMER:chipselect
	signal mm_interconnect_0_timer_s1_readdata                                : std_logic_vector(15 downto 0); -- TIMER:readdata -> mm_interconnect_0:TIMER_s1_readdata
	signal mm_interconnect_0_timer_s1_address                                 : std_logic_vector(2 downto 0);  -- mm_interconnect_0:TIMER_s1_address -> TIMER:address
	signal mm_interconnect_0_timer_s1_write                                   : std_logic;                     -- mm_interconnect_0:TIMER_s1_write -> mm_interconnect_0_timer_s1_write:in
	signal mm_interconnect_0_timer_s1_writedata                               : std_logic_vector(15 downto 0); -- mm_interconnect_0:TIMER_s1_writedata -> TIMER:writedata
	signal mm_interconnect_0_onchip_mem2_s1_chipselect                        : std_logic;                     -- mm_interconnect_0:onchip_mem2_s1_chipselect -> onchip_mem2:chipselect
	signal mm_interconnect_0_onchip_mem2_s1_readdata                          : std_logic_vector(31 downto 0); -- onchip_mem2:readdata -> mm_interconnect_0:onchip_mem2_s1_readdata
	signal mm_interconnect_0_onchip_mem2_s1_address                           : std_logic_vector(15 downto 0); -- mm_interconnect_0:onchip_mem2_s1_address -> onchip_mem2:address
	signal mm_interconnect_0_onchip_mem2_s1_byteenable                        : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_mem2_s1_byteenable -> onchip_mem2:byteenable
	signal mm_interconnect_0_onchip_mem2_s1_write                             : std_logic;                     -- mm_interconnect_0:onchip_mem2_s1_write -> onchip_mem2:write
	signal mm_interconnect_0_onchip_mem2_s1_writedata                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_mem2_s1_writedata -> onchip_mem2:writedata
	signal mm_interconnect_0_onchip_mem2_s1_clken                             : std_logic;                     -- mm_interconnect_0:onchip_mem2_s1_clken -> onchip_mem2:clken
	signal mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_readdata   : std_logic_vector(31 downto 0); -- PIXEL_BUFFER_DMA:slave_readdata -> mm_interconnect_0:PIXEL_BUFFER_DMA_avalon_control_slave_readdata
	signal mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_address    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:PIXEL_BUFFER_DMA_avalon_control_slave_address -> PIXEL_BUFFER_DMA:slave_address
	signal mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_read       : std_logic;                     -- mm_interconnect_0:PIXEL_BUFFER_DMA_avalon_control_slave_read -> PIXEL_BUFFER_DMA:slave_read
	signal mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_byteenable : std_logic_vector(3 downto 0);  -- mm_interconnect_0:PIXEL_BUFFER_DMA_avalon_control_slave_byteenable -> PIXEL_BUFFER_DMA:slave_byteenable
	signal mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_write      : std_logic;                     -- mm_interconnect_0:PIXEL_BUFFER_DMA_avalon_control_slave_write -> PIXEL_BUFFER_DMA:slave_write
	signal mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_writedata  : std_logic_vector(31 downto 0); -- mm_interconnect_0:PIXEL_BUFFER_DMA_avalon_control_slave_writedata -> PIXEL_BUFFER_DMA:slave_writedata
	signal mm_interconnect_0_nios2_vga_debug_mem_slave_readdata               : std_logic_vector(31 downto 0); -- NIOS2_VGA:debug_mem_slave_readdata -> mm_interconnect_0:NIOS2_VGA_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_vga_debug_mem_slave_waitrequest            : std_logic;                     -- NIOS2_VGA:debug_mem_slave_waitrequest -> mm_interconnect_0:NIOS2_VGA_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_vga_debug_mem_slave_debugaccess            : std_logic;                     -- mm_interconnect_0:NIOS2_VGA_debug_mem_slave_debugaccess -> NIOS2_VGA:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_vga_debug_mem_slave_address                : std_logic_vector(8 downto 0);  -- mm_interconnect_0:NIOS2_VGA_debug_mem_slave_address -> NIOS2_VGA:debug_mem_slave_address
	signal mm_interconnect_0_nios2_vga_debug_mem_slave_read                   : std_logic;                     -- mm_interconnect_0:NIOS2_VGA_debug_mem_slave_read -> NIOS2_VGA:debug_mem_slave_read
	signal mm_interconnect_0_nios2_vga_debug_mem_slave_byteenable             : std_logic_vector(3 downto 0);  -- mm_interconnect_0:NIOS2_VGA_debug_mem_slave_byteenable -> NIOS2_VGA:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_vga_debug_mem_slave_write                  : std_logic;                     -- mm_interconnect_0:NIOS2_VGA_debug_mem_slave_write -> NIOS2_VGA:debug_mem_slave_write
	signal mm_interconnect_0_nios2_vga_debug_mem_slave_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_0:NIOS2_VGA_debug_mem_slave_writedata -> NIOS2_VGA:debug_mem_slave_writedata
	signal mm_interconnect_0_onchip_mem3_s1_chipselect                        : std_logic;                     -- mm_interconnect_0:onchip_mem3_s1_chipselect -> onchip_mem3:chipselect
	signal mm_interconnect_0_onchip_mem3_s1_readdata                          : std_logic_vector(31 downto 0); -- onchip_mem3:readdata -> mm_interconnect_0:onchip_mem3_s1_readdata
	signal mm_interconnect_0_onchip_mem3_s1_address                           : std_logic_vector(15 downto 0); -- mm_interconnect_0:onchip_mem3_s1_address -> onchip_mem3:address
	signal mm_interconnect_0_onchip_mem3_s1_byteenable                        : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_mem3_s1_byteenable -> onchip_mem3:byteenable
	signal mm_interconnect_0_onchip_mem3_s1_write                             : std_logic;                     -- mm_interconnect_0:onchip_mem3_s1_write -> onchip_mem3:write
	signal mm_interconnect_0_onchip_mem3_s1_writedata                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_mem3_s1_writedata -> onchip_mem3:writedata
	signal mm_interconnect_0_onchip_mem3_s1_clken                             : std_logic;                     -- mm_interconnect_0:onchip_mem3_s1_clken -> onchip_mem3:clken
	signal nios2_nn_irq_irq                                                   : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> NIOS2_NN:irq
	signal nios2_vga_irq_irq                                                  : std_logic_vector(31 downto 0); -- irq_mapper_001:sender_irq -> NIOS2_VGA:irq
	signal irq_mapper_receiver1_irq                                           : std_logic;                     -- JTAG_UART:av_irq -> [irq_mapper:receiver1_irq, irq_mapper_001:receiver1_irq]
	signal irq_mapper_receiver0_irq                                           : std_logic;                     -- TIMER:irq -> [irq_mapper:receiver0_irq, irq_mapper_001:receiver0_irq]
	signal scaler_avalon_scaler_source_valid                                  : std_logic;                     -- SCALER:stream_out_valid -> avalon_st_adapter:in_0_valid
	signal scaler_avalon_scaler_source_data                                   : std_logic_vector(29 downto 0); -- SCALER:stream_out_data -> avalon_st_adapter:in_0_data
	signal scaler_avalon_scaler_source_ready                                  : std_logic;                     -- avalon_st_adapter:in_0_ready -> SCALER:stream_out_ready
	signal scaler_avalon_scaler_source_channel                                : std_logic_vector(1 downto 0);  -- SCALER:stream_out_channel -> avalon_st_adapter:in_0_channel
	signal scaler_avalon_scaler_source_startofpacket                          : std_logic;                     -- SCALER:stream_out_startofpacket -> avalon_st_adapter:in_0_startofpacket
	signal scaler_avalon_scaler_source_endofpacket                            : std_logic;                     -- SCALER:stream_out_endofpacket -> avalon_st_adapter:in_0_endofpacket
	signal avalon_st_adapter_out_0_valid                                      : std_logic;                     -- avalon_st_adapter:out_0_valid -> DUAL_CLOCK_FIFO:stream_in_valid
	signal avalon_st_adapter_out_0_data                                       : std_logic_vector(29 downto 0); -- avalon_st_adapter:out_0_data -> DUAL_CLOCK_FIFO:stream_in_data
	signal avalon_st_adapter_out_0_ready                                      : std_logic;                     -- DUAL_CLOCK_FIFO:stream_in_ready -> avalon_st_adapter:out_0_ready
	signal avalon_st_adapter_out_0_startofpacket                              : std_logic;                     -- avalon_st_adapter:out_0_startofpacket -> DUAL_CLOCK_FIFO:stream_in_startofpacket
	signal avalon_st_adapter_out_0_endofpacket                                : std_logic;                     -- avalon_st_adapter:out_0_endofpacket -> DUAL_CLOCK_FIFO:stream_in_endofpacket
	signal rst_controller_reset_out_reset                                     : std_logic;                     -- rst_controller:reset_out -> [DUAL_CLOCK_FIFO:reset_stream_in, PIXEL_BUFFER_DMA:reset, RGB_RESAMPLER:reset, SCALER:reset, avalon_st_adapter:in_rst_0_reset, irq_mapper:reset, irq_mapper_001:reset, mm_interconnect_0:PIXEL_BUFFER_DMA_reset_reset_bridge_in_reset_reset, onchip_mem2:reset, onchip_mem3:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                                 : std_logic;                     -- rst_controller:reset_req -> [NIOS2_NN:reset_req, NIOS2_VGA:reset_req, onchip_mem2:reset_req, onchip_mem3:reset_req, rst_translator:reset_req_in]
	signal nios2_nn_debug_reset_request_reset                                 : std_logic;                     -- NIOS2_NN:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	signal nios2_vga_debug_reset_request_reset                                : std_logic;                     -- NIOS2_VGA:debug_reset_request -> [rst_controller:reset_in2, rst_controller_001:reset_in2, rst_controller_002:reset_in2]
	signal rst_controller_001_reset_out_reset                                 : std_logic;                     -- rst_controller_001:reset_out -> [DUAL_CLOCK_FIFO:reset_stream_out, VGA:reset]
	signal rst_controller_002_reset_out_reset                                 : std_logic;                     -- rst_controller_002:reset_out -> PLL:rst
	signal reset_reset_n_ports_inv                                            : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0]
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv       : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> JTAG_UART:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv      : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> JTAG_UART:av_write_n
	signal mm_interconnect_0_sdram_vga_s1_read_ports_inv                      : std_logic;                     -- mm_interconnect_0_sdram_vga_s1_read:inv -> SDRAM_VGA:az_rd_n
	signal mm_interconnect_0_sdram_vga_s1_byteenable_ports_inv                : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_vga_s1_byteenable:inv -> SDRAM_VGA:az_be_n
	signal mm_interconnect_0_sdram_vga_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_sdram_vga_s1_write:inv -> SDRAM_VGA:az_wr_n
	signal mm_interconnect_0_timer_s1_write_ports_inv                         : std_logic;                     -- mm_interconnect_0_timer_s1_write:inv -> TIMER:write_n
	signal rst_controller_reset_out_reset_ports_inv                           : std_logic;                     -- rst_controller_reset_out_reset:inv -> [JTAG_UART:rst_n, NIOS2_NN:reset_n, NIOS2_VGA:reset_n, SDRAM_VGA:reset_n, SYSTEM_ID_1:reset_n, TIMER:reset_n, uart_0:reset_n]

begin

	dual_clock_fifo : component Sistema_Epy_DUAL_CLOCK_FIFO
		port map (
			clk_stream_in            => pll_outclk0_clk,                                       --         clock_stream_in.clk
			reset_stream_in          => rst_controller_reset_out_reset,                        --         reset_stream_in.reset
			clk_stream_out           => pll_outclk1_clk,                                       --        clock_stream_out.clk
			reset_stream_out         => rst_controller_001_reset_out_reset,                    --        reset_stream_out.reset
			stream_in_ready          => avalon_st_adapter_out_0_ready,                         --   avalon_dc_buffer_sink.ready
			stream_in_startofpacket  => avalon_st_adapter_out_0_startofpacket,                 --                        .startofpacket
			stream_in_endofpacket    => avalon_st_adapter_out_0_endofpacket,                   --                        .endofpacket
			stream_in_valid          => avalon_st_adapter_out_0_valid,                         --                        .valid
			stream_in_data           => avalon_st_adapter_out_0_data,                          --                        .data
			stream_out_ready         => dual_clock_fifo_avalon_dc_buffer_source_ready,         -- avalon_dc_buffer_source.ready
			stream_out_startofpacket => dual_clock_fifo_avalon_dc_buffer_source_startofpacket, --                        .startofpacket
			stream_out_endofpacket   => dual_clock_fifo_avalon_dc_buffer_source_endofpacket,   --                        .endofpacket
			stream_out_valid         => dual_clock_fifo_avalon_dc_buffer_source_valid,         --                        .valid
			stream_out_data          => dual_clock_fifo_avalon_dc_buffer_source_data           --                        .data
		);

	jtag_uart : component Sistema_Epy_JTAG_UART
		port map (
			clk            => pll_outclk0_clk,                                               --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver1_irq                                       --               irq.irq
		);

	nios2_nn : component Sistema_Epy_NIOS2_NN
		port map (
			clk                                 => pll_outclk0_clk,                                        --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,               --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                     --                          .reset_req
			d_address                           => nios2_nn_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_nn_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_nn_data_master_read,                              --                          .read
			d_readdata                          => nios2_nn_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_nn_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_nn_data_master_write,                             --                          .write
			d_writedata                         => nios2_nn_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios2_nn_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_nn_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_nn_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_nn_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_nn_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => nios2_nn_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_nn_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_nn_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_nn_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_nn_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_nn_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_nn_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_nn_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_nn_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_nn_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                    -- custom_instruction_master.readra
		);

	nios2_vga : component Sistema_Epy_NIOS2_VGA
		port map (
			clk                                 => pll_outclk0_clk,                                         --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,                --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                      --                          .reset_req
			d_address                           => nios2_vga_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_vga_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_vga_data_master_read,                              --                          .read
			d_readdata                          => nios2_vga_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_vga_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_vga_data_master_write,                             --                          .write
			d_writedata                         => nios2_vga_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => nios2_vga_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => nios2_vga_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_vga_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_vga_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_vga_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_vga_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => nios2_vga_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => nios2_vga_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_vga_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_vga_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_vga_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_vga_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_vga_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_vga_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_vga_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_vga_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_vga_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                     -- custom_instruction_master.readra
		);

	pixel_buffer_dma : component Sistema_Epy_PIXEL_BUFFER_DMA
		port map (
			clk                  => pll_outclk0_clk,                                                    --                     clk.clk
			reset                => rst_controller_reset_out_reset,                                     --                   reset.reset
			master_readdatavalid => pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid,             -- avalon_pixel_dma_master.readdatavalid
			master_waitrequest   => pixel_buffer_dma_avalon_pixel_dma_master_waitrequest,               --                        .waitrequest
			master_address       => pixel_buffer_dma_avalon_pixel_dma_master_address,                   --                        .address
			master_arbiterlock   => pixel_buffer_dma_avalon_pixel_dma_master_lock,                      --                        .lock
			master_read          => pixel_buffer_dma_avalon_pixel_dma_master_read,                      --                        .read
			master_readdata      => pixel_buffer_dma_avalon_pixel_dma_master_readdata,                  --                        .readdata
			slave_address        => mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_address,    --    avalon_control_slave.address
			slave_byteenable     => mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_byteenable, --                        .byteenable
			slave_read           => mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_read,       --                        .read
			slave_write          => mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_write,      --                        .write
			slave_writedata      => mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_writedata,  --                        .writedata
			slave_readdata       => mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_readdata,   --                        .readdata
			stream_ready         => pixel_buffer_dma_avalon_pixel_source_ready,                         --     avalon_pixel_source.ready
			stream_startofpacket => pixel_buffer_dma_avalon_pixel_source_startofpacket,                 --                        .startofpacket
			stream_endofpacket   => pixel_buffer_dma_avalon_pixel_source_endofpacket,                   --                        .endofpacket
			stream_valid         => pixel_buffer_dma_avalon_pixel_source_valid,                         --                        .valid
			stream_data          => pixel_buffer_dma_avalon_pixel_source_data                           --                        .data
		);

	pll : component Sistema_Epy_PLL
		port map (
			refclk   => clk_clk,                            --  refclk.clk
			rst      => rst_controller_002_reset_out_reset, --   reset.reset
			outclk_0 => pll_outclk0_clk,                    -- outclk0.clk
			outclk_1 => pll_outclk1_clk,                    -- outclk1.clk
			outclk_2 => clk_sdram_clk,                      -- outclk2.clk
			locked   => open                                -- (terminated)
		);

	rgb_resampler : component Sistema_Epy_RGB_RESAMPLER
		port map (
			clk                      => pll_outclk0_clk,                                    --               clk.clk
			reset                    => rst_controller_reset_out_reset,                     --             reset.reset
			stream_in_startofpacket  => pixel_buffer_dma_avalon_pixel_source_startofpacket, --   avalon_rgb_sink.startofpacket
			stream_in_endofpacket    => pixel_buffer_dma_avalon_pixel_source_endofpacket,   --                  .endofpacket
			stream_in_valid          => pixel_buffer_dma_avalon_pixel_source_valid,         --                  .valid
			stream_in_ready          => pixel_buffer_dma_avalon_pixel_source_ready,         --                  .ready
			stream_in_data           => pixel_buffer_dma_avalon_pixel_source_data,          --                  .data
			stream_out_ready         => rgb_resampler_avalon_rgb_source_ready,              -- avalon_rgb_source.ready
			stream_out_startofpacket => rgb_resampler_avalon_rgb_source_startofpacket,      --                  .startofpacket
			stream_out_endofpacket   => rgb_resampler_avalon_rgb_source_endofpacket,        --                  .endofpacket
			stream_out_valid         => rgb_resampler_avalon_rgb_source_valid,              --                  .valid
			stream_out_data          => rgb_resampler_avalon_rgb_source_data                --                  .data
		);

	scaler : component Sistema_Epy_SCALER
		port map (
			clk                      => pll_outclk0_clk,                               --                  clk.clk
			reset                    => rst_controller_reset_out_reset,                --                reset.reset
			stream_in_startofpacket  => rgb_resampler_avalon_rgb_source_startofpacket, --   avalon_scaler_sink.startofpacket
			stream_in_endofpacket    => rgb_resampler_avalon_rgb_source_endofpacket,   --                     .endofpacket
			stream_in_valid          => rgb_resampler_avalon_rgb_source_valid,         --                     .valid
			stream_in_ready          => rgb_resampler_avalon_rgb_source_ready,         --                     .ready
			stream_in_data           => rgb_resampler_avalon_rgb_source_data,          --                     .data
			stream_out_ready         => scaler_avalon_scaler_source_ready,             -- avalon_scaler_source.ready
			stream_out_startofpacket => scaler_avalon_scaler_source_startofpacket,     --                     .startofpacket
			stream_out_endofpacket   => scaler_avalon_scaler_source_endofpacket,       --                     .endofpacket
			stream_out_valid         => scaler_avalon_scaler_source_valid,             --                     .valid
			stream_out_data          => scaler_avalon_scaler_source_data,              --                     .data
			stream_out_channel       => scaler_avalon_scaler_source_channel            --                     .channel
		);

	sdram_vga : component Sistema_Epy_SDRAM_VGA
		port map (
			clk            => pll_outclk0_clk,                                     --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,            -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_vga_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_vga_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_vga_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_vga_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_vga_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_vga_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_vga_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_vga_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_vga_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_wire_addr,                                     --  wire.export
			zs_ba          => sdram_wire_ba,                                       --      .export
			zs_cas_n       => sdram_wire_cas_n,                                    --      .export
			zs_cke         => sdram_wire_cke,                                      --      .export
			zs_cs_n        => sdram_wire_cs_n,                                     --      .export
			zs_dq          => sdram_wire_dq,                                       --      .export
			zs_dqm         => sdram_wire_dqm,                                      --      .export
			zs_ras_n       => sdram_wire_ras_n,                                    --      .export
			zs_we_n        => sdram_wire_we_n                                      --      .export
		);

	system_id_1 : component Sistema_Epy_SYSTEM_ID_1
		port map (
			clock    => pll_outclk0_clk,                                        --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,               --         reset.reset_n
			readdata => mm_interconnect_0_system_id_1_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_system_id_1_control_slave_address(0)  --              .address
		);

	timer : component Sistema_Epy_TIMER
		port map (
			clk        => pll_outclk0_clk,                            --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   -- reset.reset_n
			address    => mm_interconnect_0_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver0_irq                    --   irq.irq
		);

	vga : component Sistema_Epy_VGA
		port map (
			clk           => pll_outclk1_clk,                                       --                clk.clk
			reset         => rst_controller_001_reset_out_reset,                    --              reset.reset
			data          => dual_clock_fifo_avalon_dc_buffer_source_data,          --    avalon_vga_sink.data
			startofpacket => dual_clock_fifo_avalon_dc_buffer_source_startofpacket, --                   .startofpacket
			endofpacket   => dual_clock_fifo_avalon_dc_buffer_source_endofpacket,   --                   .endofpacket
			valid         => dual_clock_fifo_avalon_dc_buffer_source_valid,         --                   .valid
			ready         => dual_clock_fifo_avalon_dc_buffer_source_ready,         --                   .ready
			VGA_CLK       => vga_external_interface_CLK,                            -- external_interface.export
			VGA_HS        => vga_external_interface_HS,                             --                   .export
			VGA_VS        => vga_external_interface_VS,                             --                   .export
			VGA_BLANK     => vga_external_interface_BLANK,                          --                   .export
			VGA_SYNC      => vga_external_interface_SYNC,                           --                   .export
			VGA_R         => vga_external_interface_R,                              --                   .export
			VGA_G         => vga_external_interface_G,                              --                   .export
			VGA_B         => vga_external_interface_B                               --                   .export
		);

	onchip_mem2 : component Sistema_Epy_onchip_mem2
		port map (
			clk        => pll_outclk0_clk,                             --   clk1.clk
			address    => mm_interconnect_0_onchip_mem2_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_mem2_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_mem2_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_mem2_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_mem2_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_mem2_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_mem2_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,              -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,          --       .reset_req
			freeze     => '0'                                          -- (terminated)
		);

	onchip_mem3 : component Sistema_Epy_onchip_mem3
		port map (
			clk        => pll_outclk0_clk,                             --   clk1.clk
			address    => mm_interconnect_0_onchip_mem3_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_mem3_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_mem3_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_mem3_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_mem3_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_mem3_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_mem3_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,              -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,          --       .reset_req
			freeze     => '0'                                          -- (terminated)
		);

	uart_0 : component Sistema_Epy_uart_0
		port map (
			clk           => pll_outclk0_clk,                          --                 clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address       => open,                                     --                  s1.address
			begintransfer => open,                                     --                    .begintransfer
			chipselect    => open,                                     --                    .chipselect
			read_n        => open,                                     --                    .read_n
			write_n       => open,                                     --                    .write_n
			writedata     => open,                                     --                    .writedata
			readdata      => open,                                     --                    .readdata
			rxd           => uart_rxd,                                 -- external_connection.export
			txd           => uart_txd,                                 --                    .export
			irq           => open                                      --                 irq.irq
		);

	mm_interconnect_0 : component Sistema_Epy_mm_interconnect_0
		port map (
			PLL_outclk0_clk                                        => pll_outclk0_clk,                                                    --                                  PLL_outclk0.clk
			PIXEL_BUFFER_DMA_reset_reset_bridge_in_reset_reset     => rst_controller_reset_out_reset,                                     -- PIXEL_BUFFER_DMA_reset_reset_bridge_in_reset.reset
			NIOS2_NN_data_master_address                           => nios2_nn_data_master_address,                                       --                         NIOS2_NN_data_master.address
			NIOS2_NN_data_master_waitrequest                       => nios2_nn_data_master_waitrequest,                                   --                                             .waitrequest
			NIOS2_NN_data_master_byteenable                        => nios2_nn_data_master_byteenable,                                    --                                             .byteenable
			NIOS2_NN_data_master_read                              => nios2_nn_data_master_read,                                          --                                             .read
			NIOS2_NN_data_master_readdata                          => nios2_nn_data_master_readdata,                                      --                                             .readdata
			NIOS2_NN_data_master_write                             => nios2_nn_data_master_write,                                         --                                             .write
			NIOS2_NN_data_master_writedata                         => nios2_nn_data_master_writedata,                                     --                                             .writedata
			NIOS2_NN_data_master_debugaccess                       => nios2_nn_data_master_debugaccess,                                   --                                             .debugaccess
			NIOS2_NN_instruction_master_address                    => nios2_nn_instruction_master_address,                                --                  NIOS2_NN_instruction_master.address
			NIOS2_NN_instruction_master_waitrequest                => nios2_nn_instruction_master_waitrequest,                            --                                             .waitrequest
			NIOS2_NN_instruction_master_read                       => nios2_nn_instruction_master_read,                                   --                                             .read
			NIOS2_NN_instruction_master_readdata                   => nios2_nn_instruction_master_readdata,                               --                                             .readdata
			NIOS2_VGA_data_master_address                          => nios2_vga_data_master_address,                                      --                        NIOS2_VGA_data_master.address
			NIOS2_VGA_data_master_waitrequest                      => nios2_vga_data_master_waitrequest,                                  --                                             .waitrequest
			NIOS2_VGA_data_master_byteenable                       => nios2_vga_data_master_byteenable,                                   --                                             .byteenable
			NIOS2_VGA_data_master_read                             => nios2_vga_data_master_read,                                         --                                             .read
			NIOS2_VGA_data_master_readdata                         => nios2_vga_data_master_readdata,                                     --                                             .readdata
			NIOS2_VGA_data_master_readdatavalid                    => nios2_vga_data_master_readdatavalid,                                --                                             .readdatavalid
			NIOS2_VGA_data_master_write                            => nios2_vga_data_master_write,                                        --                                             .write
			NIOS2_VGA_data_master_writedata                        => nios2_vga_data_master_writedata,                                    --                                             .writedata
			NIOS2_VGA_data_master_debugaccess                      => nios2_vga_data_master_debugaccess,                                  --                                             .debugaccess
			NIOS2_VGA_instruction_master_address                   => nios2_vga_instruction_master_address,                               --                 NIOS2_VGA_instruction_master.address
			NIOS2_VGA_instruction_master_waitrequest               => nios2_vga_instruction_master_waitrequest,                           --                                             .waitrequest
			NIOS2_VGA_instruction_master_read                      => nios2_vga_instruction_master_read,                                  --                                             .read
			NIOS2_VGA_instruction_master_readdata                  => nios2_vga_instruction_master_readdata,                              --                                             .readdata
			NIOS2_VGA_instruction_master_readdatavalid             => nios2_vga_instruction_master_readdatavalid,                         --                                             .readdatavalid
			PIXEL_BUFFER_DMA_avalon_pixel_dma_master_address       => pixel_buffer_dma_avalon_pixel_dma_master_address,                   --     PIXEL_BUFFER_DMA_avalon_pixel_dma_master.address
			PIXEL_BUFFER_DMA_avalon_pixel_dma_master_waitrequest   => pixel_buffer_dma_avalon_pixel_dma_master_waitrequest,               --                                             .waitrequest
			PIXEL_BUFFER_DMA_avalon_pixel_dma_master_read          => pixel_buffer_dma_avalon_pixel_dma_master_read,                      --                                             .read
			PIXEL_BUFFER_DMA_avalon_pixel_dma_master_readdata      => pixel_buffer_dma_avalon_pixel_dma_master_readdata,                  --                                             .readdata
			PIXEL_BUFFER_DMA_avalon_pixel_dma_master_readdatavalid => pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid,             --                                             .readdatavalid
			PIXEL_BUFFER_DMA_avalon_pixel_dma_master_lock          => pixel_buffer_dma_avalon_pixel_dma_master_lock,                      --                                             .lock
			JTAG_UART_avalon_jtag_slave_address                    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,              --                  JTAG_UART_avalon_jtag_slave.address
			JTAG_UART_avalon_jtag_slave_write                      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,                --                                             .write
			JTAG_UART_avalon_jtag_slave_read                       => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,                 --                                             .read
			JTAG_UART_avalon_jtag_slave_readdata                   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,             --                                             .readdata
			JTAG_UART_avalon_jtag_slave_writedata                  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,            --                                             .writedata
			JTAG_UART_avalon_jtag_slave_waitrequest                => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,          --                                             .waitrequest
			JTAG_UART_avalon_jtag_slave_chipselect                 => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,           --                                             .chipselect
			NIOS2_NN_debug_mem_slave_address                       => mm_interconnect_0_nios2_nn_debug_mem_slave_address,                 --                     NIOS2_NN_debug_mem_slave.address
			NIOS2_NN_debug_mem_slave_write                         => mm_interconnect_0_nios2_nn_debug_mem_slave_write,                   --                                             .write
			NIOS2_NN_debug_mem_slave_read                          => mm_interconnect_0_nios2_nn_debug_mem_slave_read,                    --                                             .read
			NIOS2_NN_debug_mem_slave_readdata                      => mm_interconnect_0_nios2_nn_debug_mem_slave_readdata,                --                                             .readdata
			NIOS2_NN_debug_mem_slave_writedata                     => mm_interconnect_0_nios2_nn_debug_mem_slave_writedata,               --                                             .writedata
			NIOS2_NN_debug_mem_slave_byteenable                    => mm_interconnect_0_nios2_nn_debug_mem_slave_byteenable,              --                                             .byteenable
			NIOS2_NN_debug_mem_slave_waitrequest                   => mm_interconnect_0_nios2_nn_debug_mem_slave_waitrequest,             --                                             .waitrequest
			NIOS2_NN_debug_mem_slave_debugaccess                   => mm_interconnect_0_nios2_nn_debug_mem_slave_debugaccess,             --                                             .debugaccess
			NIOS2_VGA_debug_mem_slave_address                      => mm_interconnect_0_nios2_vga_debug_mem_slave_address,                --                    NIOS2_VGA_debug_mem_slave.address
			NIOS2_VGA_debug_mem_slave_write                        => mm_interconnect_0_nios2_vga_debug_mem_slave_write,                  --                                             .write
			NIOS2_VGA_debug_mem_slave_read                         => mm_interconnect_0_nios2_vga_debug_mem_slave_read,                   --                                             .read
			NIOS2_VGA_debug_mem_slave_readdata                     => mm_interconnect_0_nios2_vga_debug_mem_slave_readdata,               --                                             .readdata
			NIOS2_VGA_debug_mem_slave_writedata                    => mm_interconnect_0_nios2_vga_debug_mem_slave_writedata,              --                                             .writedata
			NIOS2_VGA_debug_mem_slave_byteenable                   => mm_interconnect_0_nios2_vga_debug_mem_slave_byteenable,             --                                             .byteenable
			NIOS2_VGA_debug_mem_slave_waitrequest                  => mm_interconnect_0_nios2_vga_debug_mem_slave_waitrequest,            --                                             .waitrequest
			NIOS2_VGA_debug_mem_slave_debugaccess                  => mm_interconnect_0_nios2_vga_debug_mem_slave_debugaccess,            --                                             .debugaccess
			onchip_mem2_s1_address                                 => mm_interconnect_0_onchip_mem2_s1_address,                           --                               onchip_mem2_s1.address
			onchip_mem2_s1_write                                   => mm_interconnect_0_onchip_mem2_s1_write,                             --                                             .write
			onchip_mem2_s1_readdata                                => mm_interconnect_0_onchip_mem2_s1_readdata,                          --                                             .readdata
			onchip_mem2_s1_writedata                               => mm_interconnect_0_onchip_mem2_s1_writedata,                         --                                             .writedata
			onchip_mem2_s1_byteenable                              => mm_interconnect_0_onchip_mem2_s1_byteenable,                        --                                             .byteenable
			onchip_mem2_s1_chipselect                              => mm_interconnect_0_onchip_mem2_s1_chipselect,                        --                                             .chipselect
			onchip_mem2_s1_clken                                   => mm_interconnect_0_onchip_mem2_s1_clken,                             --                                             .clken
			onchip_mem3_s1_address                                 => mm_interconnect_0_onchip_mem3_s1_address,                           --                               onchip_mem3_s1.address
			onchip_mem3_s1_write                                   => mm_interconnect_0_onchip_mem3_s1_write,                             --                                             .write
			onchip_mem3_s1_readdata                                => mm_interconnect_0_onchip_mem3_s1_readdata,                          --                                             .readdata
			onchip_mem3_s1_writedata                               => mm_interconnect_0_onchip_mem3_s1_writedata,                         --                                             .writedata
			onchip_mem3_s1_byteenable                              => mm_interconnect_0_onchip_mem3_s1_byteenable,                        --                                             .byteenable
			onchip_mem3_s1_chipselect                              => mm_interconnect_0_onchip_mem3_s1_chipselect,                        --                                             .chipselect
			onchip_mem3_s1_clken                                   => mm_interconnect_0_onchip_mem3_s1_clken,                             --                                             .clken
			PIXEL_BUFFER_DMA_avalon_control_slave_address          => mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_address,    --        PIXEL_BUFFER_DMA_avalon_control_slave.address
			PIXEL_BUFFER_DMA_avalon_control_slave_write            => mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_write,      --                                             .write
			PIXEL_BUFFER_DMA_avalon_control_slave_read             => mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_read,       --                                             .read
			PIXEL_BUFFER_DMA_avalon_control_slave_readdata         => mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_readdata,   --                                             .readdata
			PIXEL_BUFFER_DMA_avalon_control_slave_writedata        => mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_writedata,  --                                             .writedata
			PIXEL_BUFFER_DMA_avalon_control_slave_byteenable       => mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_byteenable, --                                             .byteenable
			SDRAM_VGA_s1_address                                   => mm_interconnect_0_sdram_vga_s1_address,                             --                                 SDRAM_VGA_s1.address
			SDRAM_VGA_s1_write                                     => mm_interconnect_0_sdram_vga_s1_write,                               --                                             .write
			SDRAM_VGA_s1_read                                      => mm_interconnect_0_sdram_vga_s1_read,                                --                                             .read
			SDRAM_VGA_s1_readdata                                  => mm_interconnect_0_sdram_vga_s1_readdata,                            --                                             .readdata
			SDRAM_VGA_s1_writedata                                 => mm_interconnect_0_sdram_vga_s1_writedata,                           --                                             .writedata
			SDRAM_VGA_s1_byteenable                                => mm_interconnect_0_sdram_vga_s1_byteenable,                          --                                             .byteenable
			SDRAM_VGA_s1_readdatavalid                             => mm_interconnect_0_sdram_vga_s1_readdatavalid,                       --                                             .readdatavalid
			SDRAM_VGA_s1_waitrequest                               => mm_interconnect_0_sdram_vga_s1_waitrequest,                         --                                             .waitrequest
			SDRAM_VGA_s1_chipselect                                => mm_interconnect_0_sdram_vga_s1_chipselect,                          --                                             .chipselect
			SYSTEM_ID_1_control_slave_address                      => mm_interconnect_0_system_id_1_control_slave_address,                --                    SYSTEM_ID_1_control_slave.address
			SYSTEM_ID_1_control_slave_readdata                     => mm_interconnect_0_system_id_1_control_slave_readdata,               --                                             .readdata
			TIMER_s1_address                                       => mm_interconnect_0_timer_s1_address,                                 --                                     TIMER_s1.address
			TIMER_s1_write                                         => mm_interconnect_0_timer_s1_write,                                   --                                             .write
			TIMER_s1_readdata                                      => mm_interconnect_0_timer_s1_readdata,                                --                                             .readdata
			TIMER_s1_writedata                                     => mm_interconnect_0_timer_s1_writedata,                               --                                             .writedata
			TIMER_s1_chipselect                                    => mm_interconnect_0_timer_s1_chipselect                               --                                             .chipselect
		);

	irq_mapper : component Sistema_Epy_irq_mapper
		port map (
			clk           => pll_outclk0_clk,                --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			sender_irq    => nios2_nn_irq_irq                --    sender.irq
		);

	irq_mapper_001 : component Sistema_Epy_irq_mapper
		port map (
			clk           => pll_outclk0_clk,                --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			sender_irq    => nios2_vga_irq_irq               --    sender.irq
		);

	avalon_st_adapter : component Sistema_Epy_avalon_st_adapter
		generic map (
			inBitsPerSymbol => 10,
			inUsePackets    => 1,
			inDataWidth     => 30,
			inChannelWidth  => 2,
			inErrorWidth    => 0,
			inUseEmptyPort  => 0,
			inUseValid      => 1,
			inUseReady      => 1,
			inReadyLatency  => 0,
			outDataWidth    => 30,
			outChannelWidth => 0,
			outErrorWidth   => 0,
			outUseEmptyPort => 0,
			outUseValid     => 1,
			outUseReady     => 1,
			outReadyLatency => 0
		)
		port map (
			in_clk_0_clk        => pll_outclk0_clk,                           -- in_clk_0.clk
			in_rst_0_reset      => rst_controller_reset_out_reset,            -- in_rst_0.reset
			in_0_data           => scaler_avalon_scaler_source_data,          --     in_0.data
			in_0_valid          => scaler_avalon_scaler_source_valid,         --         .valid
			in_0_ready          => scaler_avalon_scaler_source_ready,         --         .ready
			in_0_startofpacket  => scaler_avalon_scaler_source_startofpacket, --         .startofpacket
			in_0_endofpacket    => scaler_avalon_scaler_source_endofpacket,   --         .endofpacket
			in_0_channel        => scaler_avalon_scaler_source_channel,       --         .channel
			out_0_data          => avalon_st_adapter_out_0_data,              --    out_0.data
			out_0_valid         => avalon_st_adapter_out_0_valid,             --         .valid
			out_0_ready         => avalon_st_adapter_out_0_ready,             --         .ready
			out_0_startofpacket => avalon_st_adapter_out_0_startofpacket,     --         .startofpacket
			out_0_endofpacket   => avalon_st_adapter_out_0_endofpacket        --         .endofpacket
		);

	rst_controller : component sistema_epy_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 3,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,             -- reset_in0.reset
			reset_in1      => nios2_nn_debug_reset_request_reset,  -- reset_in1.reset
			reset_in2      => nios2_vga_debug_reset_request_reset, -- reset_in2.reset
			clk            => pll_outclk0_clk,                     --       clk.clk
			reset_out      => rst_controller_reset_out_reset,      -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,  --          .reset_req
			reset_req_in0  => '0',                                 -- (terminated)
			reset_req_in1  => '0',                                 -- (terminated)
			reset_req_in2  => '0',                                 -- (terminated)
			reset_in3      => '0',                                 -- (terminated)
			reset_req_in3  => '0',                                 -- (terminated)
			reset_in4      => '0',                                 -- (terminated)
			reset_req_in4  => '0',                                 -- (terminated)
			reset_in5      => '0',                                 -- (terminated)
			reset_req_in5  => '0',                                 -- (terminated)
			reset_in6      => '0',                                 -- (terminated)
			reset_req_in6  => '0',                                 -- (terminated)
			reset_in7      => '0',                                 -- (terminated)
			reset_req_in7  => '0',                                 -- (terminated)
			reset_in8      => '0',                                 -- (terminated)
			reset_req_in8  => '0',                                 -- (terminated)
			reset_in9      => '0',                                 -- (terminated)
			reset_req_in9  => '0',                                 -- (terminated)
			reset_in10     => '0',                                 -- (terminated)
			reset_req_in10 => '0',                                 -- (terminated)
			reset_in11     => '0',                                 -- (terminated)
			reset_req_in11 => '0',                                 -- (terminated)
			reset_in12     => '0',                                 -- (terminated)
			reset_req_in12 => '0',                                 -- (terminated)
			reset_in13     => '0',                                 -- (terminated)
			reset_req_in13 => '0',                                 -- (terminated)
			reset_in14     => '0',                                 -- (terminated)
			reset_req_in14 => '0',                                 -- (terminated)
			reset_in15     => '0',                                 -- (terminated)
			reset_req_in15 => '0'                                  -- (terminated)
		);

	rst_controller_001 : component sistema_epy_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 3,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,             -- reset_in0.reset
			reset_in1      => nios2_nn_debug_reset_request_reset,  -- reset_in1.reset
			reset_in2      => nios2_vga_debug_reset_request_reset, -- reset_in2.reset
			clk            => pll_outclk1_clk,                     --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,  -- reset_out.reset
			reset_req      => open,                                -- (terminated)
			reset_req_in0  => '0',                                 -- (terminated)
			reset_req_in1  => '0',                                 -- (terminated)
			reset_req_in2  => '0',                                 -- (terminated)
			reset_in3      => '0',                                 -- (terminated)
			reset_req_in3  => '0',                                 -- (terminated)
			reset_in4      => '0',                                 -- (terminated)
			reset_req_in4  => '0',                                 -- (terminated)
			reset_in5      => '0',                                 -- (terminated)
			reset_req_in5  => '0',                                 -- (terminated)
			reset_in6      => '0',                                 -- (terminated)
			reset_req_in6  => '0',                                 -- (terminated)
			reset_in7      => '0',                                 -- (terminated)
			reset_req_in7  => '0',                                 -- (terminated)
			reset_in8      => '0',                                 -- (terminated)
			reset_req_in8  => '0',                                 -- (terminated)
			reset_in9      => '0',                                 -- (terminated)
			reset_req_in9  => '0',                                 -- (terminated)
			reset_in10     => '0',                                 -- (terminated)
			reset_req_in10 => '0',                                 -- (terminated)
			reset_in11     => '0',                                 -- (terminated)
			reset_req_in11 => '0',                                 -- (terminated)
			reset_in12     => '0',                                 -- (terminated)
			reset_req_in12 => '0',                                 -- (terminated)
			reset_in13     => '0',                                 -- (terminated)
			reset_req_in13 => '0',                                 -- (terminated)
			reset_in14     => '0',                                 -- (terminated)
			reset_req_in14 => '0',                                 -- (terminated)
			reset_in15     => '0',                                 -- (terminated)
			reset_req_in15 => '0'                                  -- (terminated)
		);

	rst_controller_002 : component sistema_epy_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 3,
			OUTPUT_RESET_SYNC_EDGES   => "none",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,             -- reset_in0.reset
			reset_in1      => nios2_nn_debug_reset_request_reset,  -- reset_in1.reset
			reset_in2      => nios2_vga_debug_reset_request_reset, -- reset_in2.reset
			clk            => open,                                --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset,  -- reset_out.reset
			reset_req      => open,                                -- (terminated)
			reset_req_in0  => '0',                                 -- (terminated)
			reset_req_in1  => '0',                                 -- (terminated)
			reset_req_in2  => '0',                                 -- (terminated)
			reset_in3      => '0',                                 -- (terminated)
			reset_req_in3  => '0',                                 -- (terminated)
			reset_in4      => '0',                                 -- (terminated)
			reset_req_in4  => '0',                                 -- (terminated)
			reset_in5      => '0',                                 -- (terminated)
			reset_req_in5  => '0',                                 -- (terminated)
			reset_in6      => '0',                                 -- (terminated)
			reset_req_in6  => '0',                                 -- (terminated)
			reset_in7      => '0',                                 -- (terminated)
			reset_req_in7  => '0',                                 -- (terminated)
			reset_in8      => '0',                                 -- (terminated)
			reset_req_in8  => '0',                                 -- (terminated)
			reset_in9      => '0',                                 -- (terminated)
			reset_req_in9  => '0',                                 -- (terminated)
			reset_in10     => '0',                                 -- (terminated)
			reset_req_in10 => '0',                                 -- (terminated)
			reset_in11     => '0',                                 -- (terminated)
			reset_req_in11 => '0',                                 -- (terminated)
			reset_in12     => '0',                                 -- (terminated)
			reset_req_in12 => '0',                                 -- (terminated)
			reset_in13     => '0',                                 -- (terminated)
			reset_req_in13 => '0',                                 -- (terminated)
			reset_in14     => '0',                                 -- (terminated)
			reset_req_in14 => '0',                                 -- (terminated)
			reset_in15     => '0',                                 -- (terminated)
			reset_req_in15 => '0'                                  -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_sdram_vga_s1_read_ports_inv <= not mm_interconnect_0_sdram_vga_s1_read;

	mm_interconnect_0_sdram_vga_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_vga_s1_byteenable;

	mm_interconnect_0_sdram_vga_s1_write_ports_inv <= not mm_interconnect_0_sdram_vga_s1_write;

	mm_interconnect_0_timer_s1_write_ports_inv <= not mm_interconnect_0_timer_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of Sistema_Epy
